`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:18:00 12/14/2017 
// Design Name: 
// Module Name:    vga_top 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
// Date: 04/04/2020
// Author: Yue (Julien) Niu
// Description: Port from NEXYS3 to NEXYS4
//////////////////////////////////////////////////////////////////////////////////
module vga_top(
	input ClkPort,
	input BtnC,
	input BtnU,
	input BtnL,
	input BtnR,

	input Sw7,
	input Sw6,
	input Sw5,
	input Sw4, 
	input Sw3, 
	input Sw2, 
	input Sw1, 
	input Sw0, // 8 switches
	
	//VGA signal
	output hSync, vSync,
	output [3:0] vgaR, vgaG, vgaB,
	
	//SSG signal 
	output An0, An1, An2, An3, An4, An5, An6, An7,
	output Ca, Cb, Cc, Cd, Ce, Cf, Cg, Dp,
	
	//output MemOE, MemWR, RamCS, 
	output QuadSpiFlashCS
	);

	// to produce divided clock
	reg [26:0]	DIV_CLK;

	assign Reset = BtnC;
	reg [7:0] Ain;
	
	wire bright;
	wire[9:0] hc, vc;
	wire[15:0] score;
	wire [6:0] ssdOut;
	wire [3:0] anode;
	wire [11:0] rgb;

	display_controller dc(.clk(ClkPort), .hSync(hSync), .vSync(vSync), .bright(bright), .hCount(hc), .vCount(vc));
	
	// use a slower clock for vga_bitchange 
	// always @(posedge ClkPort, posedge Reset) begin
	// 	if (Reset)
	// 	DIV_CLK <= 0;
    //     else
	// 	DIV_CLK <= DIV_CLK + 1'b1;
	// end

	always @(posedge ClkPort) begin
		if (Reset) begin
			Ain <= 8'b0; // Optional: reset value
		end else begin
			Ain <= {Sw7, Sw6, Sw5, Sw4, Sw3, Sw2, Sw1, Sw0};
		end
	end


	vga_bitchange vbc(.clk(ClkPort), .bright(bright), .btn_jump(BtnU), .rst(BtnC), .btn_left(BtnL), .btn_right(BtnR), .hCount(hc), .vCount(vc), .map_num(Ain), .rgb(rgb), .score(score));
	
	counter cnt(.clk(ClkPort), .displayNumber(score), .anode(anode), .ssdOut(ssdOut));
	
	assign Dp = 1;
	assign {Ca, Cb, Cc, Cd, Ce, Cf, Cg} = ssdOut[6 : 0];
    assign {An7, An6, An5, An4, An3, An2, An1, An0} = {4'b1111, anode};

	
	assign vgaR = rgb[11 : 8];
	assign vgaG = rgb[7  : 4];
	assign vgaB = rgb[3  : 0];
	
	// disable mamory ports
	//assign {MemOE, MemWR, RamCS, QuadSpiFlashCS} = 4'b1111;
	assign QuadSpiFlashCS = 1'b1;

endmodule
